module display_state(CounterX,CounterY,color,clk,clk_en,rst_n);

input clk;
input clk_en,rst_n;

output reg [7:0] CounterX,CounterY;
output reg [11:0] color;

// module vga_sin(CounterX,CounterY,color,clk,enable,reset,finished);
// module clear(CounterX,CounterY,clk,reset,enable,finished,color);
wire [7:0] CounterX_clear,CounterY_clear,CounterX_sin,CounterY_sin;
wire [11:0] color_clear, color_sin;
reg enable_clear,enable_sin,reset_clear,reset_sin;
wire finished_clear,finished_sin;


clear clear_module(
	.CounterX(CounterX_clear),
	.CounterY(CounterY_clear),
	.color(color_clear),
	.clk(clk),
	.enable(enable_clear),
	.reset(reset_clear),
	.finished(finished_clear));
	
vga_sin sin_module(
	.CounterX(CounterX_sin),
	.CounterY(CounterY_sin),
	.color(color_sin),
	.clk(clk),
	.enable(enable_sin),
	.reset(reset_sin),
	.finished(finished_sin));

parameter [1:0] clear_screen = 2'b00, draw_line = 2'b01;
reg [1:0] state,next_state;

initial begin
	state = clear_screen;
end

always @ (posedge clk)
begin
	if(rst_n == 1)
		state <= clear_screen;
	else
		state <= next_state;
end

always @ * // combinational circuit
	case(state)
		clear_screen:
		begin
			enable_clear = 1;
			enable_sin = 0;
			reset_sin = 0;

			CounterX = CounterX_clear;
			CounterY = CounterY_clear;
			color = color_clear;
			if(finished_clear == 0)
				next_state = clear_screen;
			else
				next_state = draw_line;
		end 
		draw_line:
		begin
			enable_sin = 1;
			enable_clear = 0;
			reset_clear = 0;

			CounterX = CounterX_sin;
			CounterY = CounterY_sin;
			color = color_sin;
			if(finished_sin == 0)
				next_state = draw_line;
			else
				next_state = clear_screen;
		end 
	endcase

endmodule
