module fifomapper(CounterX,CounterY,color,clk,read_clk,write_clk);

input CounterX,CounterY,color,clk,read_clk,write_clk;
//	data,
//	rdclk,
//	rdreq,
//	wrclk,
//	wrreq,
//	q,
//	rdempty,
//	wrempty,
//	wrfull);
//
//	input	[7:0]  data;
//	input	  rdclk;
//	input	  rdreq;
//	input	  wrclk;
//	input	  wrreq;
//	output	[7:0]  q;
//	output	  rdempty;
//	output	  wrempty;
//	output	  wrfull;


endmodule